----------------------------------------------------------------------------------
-- Xavier Marino & Clovis Durand
-- 
-- Create Date: 30.04.2017 13:00:22
-- Module Name: RAM - Behavioral
-- Project Name: Pmod OLEDrgb Manager
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity RAM is
    Port 
    ( 
        clk1        : in  STD_LOGIC;
        clk2        : in  STD_LOGIC;
        reset       : in  STD_LOGIC;
        w1          : in  STD_LOGIC;
        w2          : in  STD_LOGIC;
        address1    : in  STD_LOGIC_VECTOR (12 downto 0);
        address2    : in  STD_LOGIC_VECTOR (12 downto 0);
        data_in1    : in  STD_LOGIC_VECTOR (15 downto 0);
        data_in2    : in  STD_LOGIC_VECTOR (15 downto 0);
        data_out1   : out STD_LOGIC_VECTOR (15 downto 0);
        data_out2   : out STD_LOGIC_VECTOR (15 downto 0)
    );
end RAM;

architecture Behavioral of RAM is

    type   MEMORY is array (0 to 6143) of STD_LOGIC_VECTOR(15 downto 0);
    signal mem          : MEMORY := (
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"f7de",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"ef9d",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"ef7d",
                                        X"8607",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"8607",
                                        X"f7be",
                                        X"8607",
                                        X"8607",
                                        X"d6ba",
                                        X"ef7d",
                                        X"f79e",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef7d",
                                        X"f7be",
                                        X"f7be",
                                        X"ef7d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7be",
                                        X"ef9d",
                                        X"f7de",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"defb",
                                        X"defb",
                                        X"d6da",
                                        X"8607",
                                        X"8607",
                                        X"d6ba",
                                        X"ce79",
                                        X"8607",
                                        X"ce99",
                                        X"d6ba",
                                        X"d6ba",
                                        X"d6da",
                                        X"d6da",
                                        X"d6da",
                                        X"d6da",
                                        X"df1b",
                                        X"e73c",
                                        X"df1c",
                                        X"e73c",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9e",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7be",
                                        X"ef7d",
                                        X"df1b",
                                        X"e73c",
                                        X"8607",
                                        X"d6ba",
                                        X"ce99",
                                        X"d6ba",
                                        X"d6ba",
                                        X"c658",
                                        X"c658",
                                        X"ce9a",
                                        X"d6ba",
                                        X"8607",
                                        X"d6ba",
                                        X"d6ba",
                                        X"d69a",
                                        X"c618",
                                        X"c658",
                                        X"d6ba",
                                        X"ce79",
                                        X"d69a",
                                        X"ce99",
                                        X"c638",
                                        X"c638",
                                        X"c658",
                                        X"c658",
                                        X"c658",
                                        X"c658",
                                        X"ce79",
                                        X"d6ba",
                                        X"d6da",
                                        X"df1b",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"8607",
                                        X"8607",
                                        X"f7de",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7de",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"8607",
                                        X"e73c",
                                        X"e75c",
                                        X"defb",
                                        X"ce79",
                                        X"d6da",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"d6da",
                                        X"c658",
                                        X"e73c",
                                        X"e73c",
                                        X"8607",
                                        X"df1c",
                                        X"defb",
                                        X"e73c",
                                        X"ce59",
                                        X"ce79",
                                        X"defb",
                                        X"ce99",
                                        X"df1b",
                                        X"df1b",
                                        X"ce79",
                                        X"ce79",
                                        X"d69a",
                                        X"ce59",
                                        X"ce99",
                                        X"c638",
                                        X"ce79",
                                        X"ce59",
                                        X"c638",
                                        X"c638",
                                        X"ce79",
                                        X"d6ba",
                                        X"df1b",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"ef7d",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"df1c",
                                        X"f7be",
                                        X"ef7d",
                                        X"e73c",
                                        X"ef7d",
                                        X"e73c",
                                        X"d6db",
                                        X"d6ba",
                                        X"d6ba",
                                        X"ce79",
                                        X"d6ba",
                                        X"e75c",
                                        X"d6db",
                                        X"ce99",
                                        X"e75c",
                                        X"ef7d",
                                        X"d6ba",
                                        X"df1b",
                                        X"ef9d",
                                        X"e75c",
                                        X"ef7d",
                                        X"df1b",
                                        X"e75c",
                                        X"ce59",
                                        X"c638",
                                        X"df1c",
                                        X"d6ba",
                                        X"df1b",
                                        X"d6ba",
                                        X"c659",
                                        X"ce79",
                                        X"ce79",
                                        X"d6ba",
                                        X"d6da",
                                        X"c638",
                                        X"ce59",
                                        X"ce99",
                                        X"c658",
                                        X"ce79",
                                        X"ce59",
                                        X"ce79",
                                        X"ce79",
                                        X"d6ba",
                                        X"df1b",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef7d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"ef7d",
                                        X"ef7d",
                                        X"f7be",
                                        X"e75d",
                                        X"ef9d",
                                        X"f7de",
                                        X"f7de",
                                        X"e75c",
                                        X"d6ba",
                                        X"ef7d",
                                        X"df1b",
                                        X"ce99",
                                        X"ce79",
                                        X"ce99",
                                        X"d6da",
                                        X"e73c",
                                        X"e73c",
                                        X"d6da",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ce99",
                                        X"defb",
                                        X"f7de",
                                        X"ef7d",
                                        X"d69a",
                                        X"ef7d",
                                        X"e75c",
                                        X"e73c",
                                        X"d6ba",
                                        X"e73c",
                                        X"d6da",
                                        X"bdf7",
                                        X"defb",
                                        X"d6da",
                                        X"ce99",
                                        X"defb",
                                        X"d6da",
                                        X"ce79",
                                        X"ce99",
                                        X"d6ba",
                                        X"d6da",
                                        X"ce79",
                                        X"ce79",
                                        X"ce79",
                                        X"c658",
                                        X"ce99",
                                        X"ce9a",
                                        X"ce59",
                                        X"ce79",
                                        X"ce79",
                                        X"ce79",
                                        X"d69a",
                                        X"df1b",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef9e",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"e75d",
                                        X"f7be",
                                        X"ef9d",
                                        X"ce79",
                                        X"ce59",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"ef9d",
                                        X"ef9d",
                                        X"8607",
                                        X"df1b",
                                        X"f7be",
                                        X"e75c",
                                        X"d6ba",
                                        X"8607",
                                        X"ef7d",
                                        X"defb",
                                        X"d6ba",
                                        X"e75c",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"df1b",
                                        X"be17",
                                        X"d6ba",
                                        X"d6db",
                                        X"c658",
                                        X"d69a",
                                        X"defb",
                                        X"ce79",
                                        X"d6da",
                                        X"ce99",
                                        X"d6ba",
                                        X"c659",
                                        X"c658",
                                        X"ce79",
                                        X"ce79",
                                        X"ce59",
                                        X"ce79",
                                        X"c638",
                                        X"ce79",
                                        X"ce99",
                                        X"ce79",
                                        X"c658",
                                        X"ce79",
                                        X"ce9a",
                                        X"df1b",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"ef7d",
                                        X"f7be",
                                        X"e75c",
                                        X"8607",
                                        X"defb",
                                        X"d6db",
                                        X"ce9a",
                                        X"c618",
                                        X"ce79",
                                        X"e75c",
                                        X"8607",
                                        X"df1b",
                                        X"e73c",
                                        X"ef9d",
                                        X"ef9d",
                                        X"8607",
                                        X"8607",
                                        X"df1b",
                                        X"f7be",
                                        X"d6da",
                                        X"8607",
                                        X"d6da",
                                        X"e73c",
                                        X"ce79",
                                        X"8607",
                                        X"defb",
                                        X"defb",
                                        X"d6ba",
                                        X"8607",
                                        X"c638",
                                        X"ce99",
                                        X"d6da",
                                        X"ce79",
                                        X"ce79",
                                        X"d69a",
                                        X"c618",
                                        X"c658",
                                        X"ce79",
                                        X"ce99",
                                        X"ce9a",
                                        X"ce79",
                                        X"ce99",
                                        X"ce79",
                                        X"c638",
                                        X"c638",
                                        X"ce59",
                                        X"ce9a",
                                        X"ce79",
                                        X"ce59",
                                        X"c658",
                                        X"c658",
                                        X"c658",
                                        X"ce99",
                                        X"defb",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"d6ba",
                                        X"bdf7",
                                        X"ce79",
                                        X"e73c",
                                        X"e73c",
                                        X"c618",
                                        X"ce99",
                                        X"8607",
                                        X"ef7d",
                                        X"defb",
                                        X"d6da",
                                        X"e75c",
                                        X"8607",
                                        X"e73c",
                                        X"8607",
                                        X"d6db",
                                        X"defb",
                                        X"8607",
                                        X"e73c",
                                        X"df1c",
                                        X"ce59",
                                        X"8607",
                                        X"c638",
                                        X"ce59",
                                        X"c658",
                                        X"8607",
                                        X"be17",
                                        X"c618",
                                        X"c638",
                                        X"c638",
                                        X"c638",
                                        X"c638",
                                        X"be17",
                                        X"c659",
                                        X"ce99",
                                        X"ce99",
                                        X"defb",
                                        X"ce79",
                                        X"c659",
                                        X"ce79",
                                        X"c638",
                                        X"c618",
                                        X"ce99",
                                        X"c638",
                                        X"c638",
                                        X"c658",
                                        X"c638",
                                        X"ce79",
                                        X"c658",
                                        X"c638",
                                        X"ce79",
                                        X"d6ba",
                                        X"e73c",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f79e",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"255b",
                                        X"255b",
                                        X"255b",
                                        X"255b",
                                        X"255b",
                                        X"255b",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"f7de",
                                        X"f7be",
                                        X"f7be",
                                        X"8607",
                                        X"ef7d",
                                        X"8607",
                                        X"c638",
                                        X"d6ba",
                                        X"d6ba",
                                        X"be18",
                                        X"d6ba",
                                        X"e75c",
                                        X"d6ba",
                                        X"c658",
                                        X"8607",
                                        X"e75c",
                                        X"ef9d",
                                        X"df1b",
                                        X"d69a",
                                        X"8607",
                                        X"defb",
                                        X"defb",
                                        X"8607",
                                        X"d6da",
                                        X"8607",
                                        X"c658",
                                        X"ce79",
                                        X"ce99",
                                        X"8607",
                                        X"be17",
                                        X"c638",
                                        X"c658",
                                        X"8607",
                                        X"be17",
                                        X"bdf7",
                                        X"be17",
                                        X"be17",
                                        X"be17",
                                        X"be17",
                                        X"bdf7",
                                        X"c658",
                                        X"c638",
                                        X"c638",
                                        X"ce79",
                                        X"c658",
                                        X"c658",
                                        X"ce99",
                                        X"c659",
                                        X"ce79",
                                        X"ce79",
                                        X"be17",
                                        X"c638",
                                        X"c638",
                                        X"c638",
                                        X"ce79",
                                        X"c638",
                                        X"c638",
                                        X"ce79",
                                        X"ce79",
                                        X"d6ba",
                                        X"e73c",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7be",
                                        X"f7be",
                                        X"8607",
                                        X"defb",
                                        X"ce99",
                                        X"8607",
                                        X"ce59",
                                        X"e73c",
                                        X"e73c",
                                        X"c638",
                                        X"c658",
                                        X"ce99",
                                        X"d6da",
                                        X"8607",
                                        X"c638",
                                        X"d6da",
                                        X"d6da",
                                        X"defb",
                                        X"8607",
                                        X"ce59",
                                        X"ce79",
                                        X"ce79",
                                        X"8607",
                                        X"8607",
                                        X"c638",
                                        X"c638",
                                        X"be17",
                                        X"8607",
                                        X"bdf7",
                                        X"be17",
                                        X"bdf7",
                                        X"8607",
                                        X"c638",
                                        X"be17",
                                        X"be17",
                                        X"bdf7",
                                        X"bdf7",
                                        X"c638",
                                        X"be17",
                                        X"be17",
                                        X"be17",
                                        X"c658",
                                        X"ce79",
                                        X"c658",
                                        X"be17",
                                        X"be17",
                                        X"c638",
                                        X"ce79",
                                        X"ce79",
                                        X"ce79",
                                        X"c658",
                                        X"c638",
                                        X"c658",
                                        X"c638",
                                        X"c638",
                                        X"ce79",
                                        X"c658",
                                        X"c658",
                                        X"ce79",
                                        X"ce79",
                                        X"df1b",
                                        X"e73c",
                                        X"ef7d",
                                        X"ef9d",
                                        X"f79e",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"ef7d",
                                        X"8607",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"8607",
                                        X"ef7d",
                                        X"e73c",
                                        X"8607",
                                        X"ce99",
                                        X"d6da",
                                        X"df1b",
                                        X"8607",
                                        X"c618",
                                        X"defb",
                                        X"e73c",
                                        X"c658",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"c638",
                                        X"c658",
                                        X"8607",
                                        X"c618",
                                        X"be17",
                                        X"ce79",
                                        X"ce79",
                                        X"8607",
                                        X"c638",
                                        X"c658",
                                        X"c618",
                                        X"c638",
                                        X"8607",
                                        X"8607",
                                        X"8607",
                                        X"c638",
                                        X"c638",
                                        X"bdf7",
                                        X"be18",
                                        X"bdf7",
                                        X"be17",
                                        X"c618",
                                        X"be17",
                                        X"bdf7",
                                        X"bdf7",
                                        X"c618",
                                        X"c658",
                                        X"be18",
                                        X"be17",
                                        X"c638",
                                        X"c638",
                                        X"c658",
                                        X"c658",
                                        X"c658",
                                        X"c638",
                                        X"c638",
                                        X"c638",
                                        X"c638",
                                        X"c638",
                                        X"c638",
                                        X"be17",
                                        X"c638",
                                        X"ce79",
                                        X"ce79",
                                        X"ce99",
                                        X"defb",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"ef9d",
                                        X"df1b",
                                        X"e73c",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"f79e",
                                        X"ef9d",
                                        X"e73c",
                                        X"ce99",
                                        X"d6ba",
                                        X"defb",
                                        X"e73c",
                                        X"e75c",
                                        X"e73c",
                                        X"df1b",
                                        X"c659",
                                        X"d6da",
                                        X"df1b",
                                        X"ce79",
                                        X"c638",
                                        X"c658",
                                        X"c658",
                                        X"be17",
                                        X"c618",
                                        X"c618",
                                        X"be17",
                                        X"bdf7",
                                        X"c638",
                                        X"c659",
                                        X"c638",
                                        X"c638",
                                        X"be17",
                                        X"c618",
                                        X"c638",
                                        X"c638",
                                        X"be18",
                                        X"be18",
                                        X"be38",
                                        X"be18",
                                        X"be18",
                                        X"be37",
                                        X"be17",
                                        X"be38",
                                        X"be37",
                                        X"be17",
                                        X"c638",
                                        X"be17",
                                        X"be17",
                                        X"be17",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"be17",
                                        X"be18",
                                        X"be17",
                                        X"c618",
                                        X"c658",
                                        X"c638",
                                        X"c638",
                                        X"ce59",
                                        X"c658",
                                        X"c638",
                                        X"c618",
                                        X"bdf7",
                                        X"c618",
                                        X"c658",
                                        X"ce99",
                                        X"ce99",
                                        X"ce99",
                                        X"defb",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"ef9d",
                                        X"ef9d",
                                        X"df1b",
                                        X"f7be",
                                        X"f7be",
                                        X"ef9d",
                                        X"e73c",
                                        X"d6ba",
                                        X"d6da",
                                        X"df1c",
                                        X"e75c",
                                        X"e73c",
                                        X"ef7d",
                                        X"e75d",
                                        X"defb",
                                        X"ef7d",
                                        X"ce99",
                                        X"d6da",
                                        X"e75c",
                                        X"defb",
                                        X"c658",
                                        X"c658",
                                        X"bdf7",
                                        X"be17",
                                        X"be17",
                                        X"bdf7",
                                        X"bdf7",
                                        X"be17",
                                        X"bdf7",
                                        X"be17",
                                        X"c638",
                                        X"c638",
                                        X"be18",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"be17",
                                        X"c638",
                                        X"c637",
                                        X"c637",
                                        X"c678",
                                        X"ce78",
                                        X"c657",
                                        X"c657",
                                        X"c657",
                                        X"ce77",
                                        X"c658",
                                        X"c658",
                                        X"c638",
                                        X"be38",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"be17",
                                        X"c638",
                                        X"c638",
                                        X"be17",
                                        X"be17",
                                        X"c638",
                                        X"ce79",
                                        X"c618",
                                        X"be17",
                                        X"be17",
                                        X"be17",
                                        X"c658",
                                        X"ce59",
                                        X"c638",
                                        X"ce99",
                                        X"ce99",
                                        X"defb",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"ef9d",
                                        X"f7de",
                                        X"f7de",
                                        X"e75c",
                                        X"df1b",
                                        X"defb",
                                        X"df1b",
                                        X"df1b",
                                        X"d6da",
                                        X"defb",
                                        X"e75c",
                                        X"e73c",
                                        X"e73c",
                                        X"e75c",
                                        X"e75c",
                                        X"f7be",
                                        X"df1b",
                                        X"d6da",
                                        X"df1b",
                                        X"d6da",
                                        X"ce99",
                                        X"d6da",
                                        X"c659",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"be17",
                                        X"c638",
                                        X"be17",
                                        X"bdf7",
                                        X"be17",
                                        X"bdf7",
                                        X"bdf7",
                                        X"be18",
                                        X"be18",
                                        X"be18",
                                        X"be59",
                                        X"be38",
                                        X"be59",
                                        X"c69a",
                                        X"c699",
                                        X"cedb",
                                        X"d73c",
                                        X"d71c",
                                        X"d697",
                                        X"d698",
                                        X"d6b8",
                                        X"d6d8",
                                        X"ce78",
                                        X"c678",
                                        X"c678",
                                        X"be38",
                                        X"be18",
                                        X"be38",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"be38",
                                        X"c658",
                                        X"c638",
                                        X"ce99",
                                        X"be18",
                                        X"c638",
                                        X"c659",
                                        X"c638",
                                        X"c638",
                                        X"c638",
                                        X"c638",
                                        X"c618",
                                        X"c638",
                                        X"c658",
                                        X"ce99",
                                        X"ce9a",
                                        X"defb",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e75c",
                                        X"d6da",
                                        X"e75c",
                                        X"ce59",
                                        X"be17",
                                        X"df1b",
                                        X"ef9d",
                                        X"ef9d",
                                        X"e75c",
                                        X"e75c",
                                        X"e75c",
                                        X"ef7d",
                                        X"e75c",
                                        X"e75c",
                                        X"defb",
                                        X"d6da",
                                        X"d6da",
                                        X"d6ba",
                                        X"c638",
                                        X"be17",
                                        X"be17",
                                        X"bdf7",
                                        X"c638",
                                        X"c658",
                                        X"ce99",
                                        X"be17",
                                        X"c658",
                                        X"c618",
                                        X"bdf7",
                                        X"be18",
                                        X"be18",
                                        X"be39",
                                        X"be5a",
                                        X"bebb",
                                        X"c6db",
                                        X"cefd",
                                        X"cf3d",
                                        X"cefb",
                                        X"d73d",
                                        X"d73d",
                                        X"d73c",
                                        X"d697",
                                        X"d698",
                                        X"d6d9",
                                        X"ded8",
                                        X"deb7",
                                        X"ceb8",
                                        X"be59",
                                        X"be59",
                                        X"be79",
                                        X"be39",
                                        X"be18",
                                        X"be18",
                                        X"bdf7",
                                        X"be18",
                                        X"ce9a",
                                        X"ce99",
                                        X"ce79",
                                        X"ce79",
                                        X"ce59",
                                        X"c659",
                                        X"c638",
                                        X"c658",
                                        X"c638",
                                        X"be17",
                                        X"be17",
                                        X"c638",
                                        X"c638",
                                        X"ce59",
                                        X"ce99",
                                        X"ce79",
                                        X"defb",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"e75c",
                                        X"f7be",
                                        X"df1b",
                                        X"defb",
                                        X"d6ba",
                                        X"defb",
                                        X"d6da",
                                        X"ce79",
                                        X"d6da",
                                        X"e73c",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e75c",
                                        X"ef7d",
                                        X"e73c",
                                        X"df1b",
                                        X"e73c",
                                        X"df1b",
                                        X"ce99",
                                        X"ce59",
                                        X"c658",
                                        X"c618",
                                        X"c638",
                                        X"c658",
                                        X"be17",
                                        X"c638",
                                        X"c638",
                                        X"ce79",
                                        X"c659",
                                        X"bdf7",
                                        X"be18",
                                        X"be39",
                                        X"be7a",
                                        X"cefc",
                                        X"cf1d",
                                        X"cf3d",
                                        X"cefc",
                                        X"d75d",
                                        X"cf1d",
                                        X"cefb",
                                        X"d75d",
                                        X"d75d",
                                        X"d71c",
                                        X"ce99",
                                        X"d6fb",
                                        X"d6da",
                                        X"d6d9",
                                        X"df18",
                                        X"d719",
                                        X"c6da",
                                        X"be9a",
                                        X"be9a",
                                        X"be59",
                                        X"be5a",
                                        X"be39",
                                        X"be18",
                                        X"bdf8",
                                        X"be7a",
                                        X"d6fb",
                                        X"ce79",
                                        X"ce59",
                                        X"ce59",
                                        X"ce99",
                                        X"ce59",
                                        X"c638",
                                        X"c658",
                                        X"be17",
                                        X"bdf7",
                                        X"bdf7",
                                        X"be17",
                                        X"c638",
                                        X"c638",
                                        X"c658",
                                        X"ce79",
                                        X"df1b",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"f7de",
                                        X"ef7d",
                                        X"ef7d",
                                        X"f7de",
                                        X"defb",
                                        X"e0e4",
                                        X"ce79",
                                        X"e75c",
                                        X"d6da",
                                        X"c658",
                                        X"ce99",
                                        X"ce99",
                                        X"d6ba",
                                        X"d6da",
                                        X"d6da",
                                        X"ce99",
                                        X"ce99",
                                        X"c658",
                                        X"be17",
                                        X"be17",
                                        X"bdf7",
                                        X"be17",
                                        X"c659",
                                        X"ce99",
                                        X"be17",
                                        X"c638",
                                        X"ce99",
                                        X"df1b",
                                        X"df1b",
                                        X"be38",
                                        X"e0e4",
                                        X"be39",
                                        X"be7b",
                                        X"cefc",
                                        X"d73d",
                                        X"c6fd",
                                        X"c71d",
                                        X"bedc",
                                        X"e79e",
                                        X"e7be",
                                        X"cf3d",
                                        X"e79e",
                                        X"df9e",
                                        X"c6bc",
                                        X"be18",
                                        X"be39",
                                        X"c699",
                                        X"d73b",
                                        X"d71a",
                                        X"df39",
                                        X"ced9",
                                        X"beba",
                                        X"c6db",
                                        X"be9a",
                                        X"be5a",
                                        X"be39",
                                        X"be18",
                                        X"be18",
                                        X"be7a",
                                        X"d6fc",
                                        X"e73c",
                                        X"e75c",
                                        X"ce99",
                                        X"c658",
                                        X"d69a",
                                        X"c658",
                                        X"ce79",
                                        X"be17",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"be18",
                                        X"c658",
                                        X"ce79",
                                        X"ce99",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"f7de",
                                        X"f7be",
                                        X"f7de",
                                        X"e0e4",
                                        X"f7de",
                                        X"e75c",
                                        X"e73c",
                                        X"f7de",
                                        X"e0e4",
                                        X"ce79",
                                        X"ce99",
                                        X"d6da",
                                        X"ce9a",
                                        X"ce99",
                                        X"ce79",
                                        X"ce99",
                                        X"c618",
                                        X"c638",
                                        X"ce59",
                                        X"c659",
                                        X"be17",
                                        X"c638",
                                        X"be17",
                                        X"c638",
                                        X"ce79",
                                        X"d69a",
                                        X"be17",
                                        X"be17",
                                        X"d6da",
                                        X"e75c",
                                        X"ef7d",
                                        X"cedb",
                                        X"be39",
                                        X"be39",
                                        X"be5a",
                                        X"c6dc",
                                        X"d73d",
                                        X"d75d",
                                        X"c6dd",
                                        X"d75e",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"f7de",
                                        X"efde",
                                        X"d75e",
                                        X"be7b",
                                        X"be19",
                                        X"bdf9",
                                        X"bdf8",
                                        X"c6ba",
                                        X"d6fa",
                                        X"d719",
                                        X"d73b",
                                        X"cefc",
                                        X"bebb",
                                        X"be5a",
                                        X"be5a",
                                        X"be5a",
                                        X"be3a",
                                        X"be39",
                                        X"be5a",
                                        X"cedc",
                                        X"e73c",
                                        X"e75c",
                                        X"e73c",
                                        X"ce9a",
                                        X"ce79",
                                        X"ce99",
                                        X"d6da",
                                        X"c658",
                                        X"c638",
                                        X"be17",
                                        X"bdf7",
                                        X"bdf7",
                                        X"be17",
                                        X"be17",
                                        X"c638",
                                        X"c638",
                                        X"d6da",
                                        X"e75c",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef9d",
                                        X"f79e",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"ef9d",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"df1b",
                                        X"d6da",
                                        X"e0e4",
                                        X"e75c",
                                        X"c658",
                                        X"c658",
                                        X"c658",
                                        X"c658",
                                        X"c638",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"ce79",
                                        X"ce79",
                                        X"ce59",
                                        X"e0e4",
                                        X"ce99",
                                        X"ce79",
                                        X"be17",
                                        X"ce79",
                                        X"e0e4",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"cedb",
                                        X"be9a",
                                        X"e0e4",
                                        X"be3a",
                                        X"be7b",
                                        X"c6dc",
                                        X"df9e",
                                        X"e7be",
                                        X"e0e4",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"cefd",
                                        X"be3a",
                                        X"be19",
                                        X"be18",
                                        X"bdf8",
                                        X"bdf7",
                                        X"be18",
                                        X"ceba",
                                        X"d71b",
                                        X"d73b",
                                        X"cefb",
                                        X"be9b",
                                        X"be7b",
                                        X"be5b",
                                        X"be5a",
                                        X"be39",
                                        X"be39",
                                        X"be59",
                                        X"cedc",
                                        X"df3c",
                                        X"e75c",
                                        X"ef7d",
                                        X"e75c",
                                        X"df1b",
                                        X"d6ba",
                                        X"d6ba",
                                        X"ce79",
                                        X"ce79",
                                        X"c658",
                                        X"c638",
                                        X"be17",
                                        X"bdf7",
                                        X"be17",
                                        X"c638",
                                        X"ce59",
                                        X"ce79",
                                        X"df1b",
                                        X"e75c",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"e73c",
                                        X"e0e4",
                                        X"e73c",
                                        X"df1b",
                                        X"c658",
                                        X"c618",
                                        X"be17",
                                        X"e0e4",
                                        X"c658",
                                        X"c638",
                                        X"c638",
                                        X"be17",
                                        X"e0e4",
                                        X"c638",
                                        X"be18",
                                        X"e0e4",
                                        X"be17",
                                        X"c658",
                                        X"d6da",
                                        X"e75c",
                                        X"e0e4",
                                        X"ef9d",
                                        X"f7be",
                                        X"ef7d",
                                        X"d71c",
                                        X"c6bb",
                                        X"e0e4",
                                        X"be5a",
                                        X"be5a",
                                        X"c6fd",
                                        X"cf3d",
                                        X"df9e",
                                        X"e7be",
                                        X"e0e4",
                                        X"e0e4",
                                        X"efde",
                                        X"c71d",
                                        X"be19",
                                        X"bdf8",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"ceba",
                                        X"d6fa",
                                        X"ced9",
                                        X"cefa",
                                        X"be9b",
                                        X"be7b",
                                        X"be7b",
                                        X"be3a",
                                        X"be39",
                                        X"be59",
                                        X"be59",
                                        X"cedb",
                                        X"df3d",
                                        X"e75d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"d6da",
                                        X"ce79",
                                        X"ce79",
                                        X"ce79",
                                        X"d6ba",
                                        X"ce79",
                                        X"c638",
                                        X"bdf7",
                                        X"bdf7",
                                        X"be18",
                                        X"c658",
                                        X"ce79",
                                        X"ce99",
                                        X"e73c",
                                        X"e73c",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef9d",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"defb",
                                        X"defb",
                                        X"ef9d",
                                        X"f7be",
                                        X"e0e4",
                                        X"be17",
                                        X"d6ba",
                                        X"ce59",
                                        X"c658",
                                        X"c658",
                                        X"e0e4",
                                        X"ce79",
                                        X"be17",
                                        X"bdf7",
                                        X"be17",
                                        X"e0e4",
                                        X"be17",
                                        X"c638",
                                        X"c658",
                                        X"e0e4",
                                        X"e73c",
                                        X"ef9d",
                                        X"e0e4",
                                        X"f79e",
                                        X"f7be",
                                        X"f7be",
                                        X"e77d",
                                        X"c6dc",
                                        X"be5a",
                                        X"e0e4",
                                        X"be7b",
                                        X"be7b",
                                        X"c71d",
                                        X"d77e",
                                        X"cf5e",
                                        X"c73d",
                                        X"c71e",
                                        X"d77e",
                                        X"e0e4",
                                        X"be7a",
                                        X"bdf8",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"ce99",
                                        X"d71a",
                                        X"d73a",
                                        X"c6fb",
                                        X"bebb",
                                        X"bedc",
                                        X"be7b",
                                        X"be5a",
                                        X"be7b",
                                        X"be9a",
                                        X"be7a",
                                        X"cedb",
                                        X"df5d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e73c",
                                        X"ce59",
                                        X"d6da",
                                        X"d69a",
                                        X"ce79",
                                        X"ce99",
                                        X"ce79",
                                        X"c658",
                                        X"c618",
                                        X"be17",
                                        X"c638",
                                        X"ce79",
                                        X"ce79",
                                        X"d6ba",
                                        X"df1b",
                                        X"e75c",
                                        X"e75c",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7be",
                                        X"ef9d",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"f7be",
                                        X"f7bd",
                                        X"d6ba",
                                        X"defb",
                                        X"defb",
                                        X"e0e4",
                                        X"e0e4",
                                        X"c638",
                                        X"c638",
                                        X"c618",
                                        X"be17",
                                        X"c658",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"c658",
                                        X"c638",
                                        X"ce59",
                                        X"df1b",
                                        X"ef7d",
                                        X"e0e4",
                                        X"e0e4",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"ef9d",
                                        X"c6dc",
                                        X"be3a",
                                        X"e0e4",
                                        X"be9b",
                                        X"c6fc",
                                        X"cf3d",
                                        X"cf5e",
                                        X"d75e",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"d6fb",
                                        X"c659",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"c6ba",
                                        X"d75c",
                                        X"df7c",
                                        X"cf3b",
                                        X"bebb",
                                        X"bebc",
                                        X"be7a",
                                        X"be5a",
                                        X"be9b",
                                        X"c6ba",
                                        X"c69a",
                                        X"cedb",
                                        X"e75d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"df1b",
                                        X"ce99",
                                        X"d6ba",
                                        X"ce79",
                                        X"ce99",
                                        X"ce79",
                                        X"d6ba",
                                        X"ce99",
                                        X"be17",
                                        X"be17",
                                        X"c638",
                                        X"c638",
                                        X"ce79",
                                        X"defb",
                                        X"e73c",
                                        X"e75c",
                                        X"ef7d",
                                        X"f7be",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"ef7d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"d6ba",
                                        X"d69a",
                                        X"ce99",
                                        X"d6ba",
                                        X"ce99",
                                        X"c638",
                                        X"c618",
                                        X"c638",
                                        X"be17",
                                        X"be17",
                                        X"c638",
                                        X"be17",
                                        X"be17",
                                        X"bdf7",
                                        X"ce79",
                                        X"defb",
                                        X"e75c",
                                        X"ef7d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"efbe",
                                        X"cefc",
                                        X"be7a",
                                        X"c6db",
                                        X"d73d",
                                        X"df7e",
                                        X"d75e",
                                        X"bf1d",
                                        X"cf5e",
                                        X"d75d",
                                        X"d75d",
                                        X"cf3c",
                                        X"cefa",
                                        X"c69a",
                                        X"be3a",
                                        X"be19",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"c6db",
                                        X"df7b",
                                        X"df7b",
                                        X"d73c",
                                        X"c6fd",
                                        X"c6dd",
                                        X"be9c",
                                        X"be7b",
                                        X"be7a",
                                        X"be7a",
                                        X"be7a",
                                        X"cedc",
                                        X"e75d",
                                        X"ef9d",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"e73c",
                                        X"d6da",
                                        X"d6da",
                                        X"d6ba",
                                        X"ce79",
                                        X"ce79",
                                        X"ce9a",
                                        X"d69a",
                                        X"ce79",
                                        X"c658",
                                        X"c638",
                                        X"c618",
                                        X"c659",
                                        X"ce79",
                                        X"defb",
                                        X"e75c",
                                        X"ef7d",
                                        X"f7be",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"e73c",
                                        X"ef9d",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"e73c",
                                        X"e73c",
                                        X"d6da",
                                        X"ce79",
                                        X"ce79",
                                        X"c638",
                                        X"c618",
                                        X"c659",
                                        X"c638",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"be17",
                                        X"c638",
                                        X"d6da",
                                        X"e73c",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"efbe",
                                        X"d73d",
                                        X"c6fc",
                                        X"d71c",
                                        X"df5d",
                                        X"df9e",
                                        X"d77e",
                                        X"c73e",
                                        X"c75e",
                                        X"d75e",
                                        X"cf3d",
                                        X"cf3c",
                                        X"cf1c",
                                        X"c6bb",
                                        X"be9c",
                                        X"be5b",
                                        X"bdf8",
                                        X"bdf7",
                                        X"bdf7",
                                        X"bdf7",
                                        X"c659",
                                        X"d71b",
                                        X"df7a",
                                        X"d75a",
                                        X"bedc",
                                        X"bedc",
                                        X"bedd",
                                        X"be9c",
                                        X"bebc",
                                        X"be9b",
                                        X"be7a",
                                        X"be7a",
                                        X"d6fc",
                                        X"ef7d",
                                        X"f7be",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"e75c",
                                        X"df1b",
                                        X"d6da",
                                        X"d6ba",
                                        X"ce99",
                                        X"ce79",
                                        X"ce99",
                                        X"d6ba",
                                        X"d6ba",
                                        X"d69a",
                                        X"c659",
                                        X"ce79",
                                        X"ce79",
                                        X"c658",
                                        X"defb",
                                        X"e73c",
                                        X"ef7d",
                                        X"f7be",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"f7de",
                                        X"f7be",
                                        X"e73c",
                                        X"e0e4",
                                        X"d6da",
                                        X"d6da",
                                        X"d6da",
                                        X"ce59",
                                        X"e0e4",
                                        X"bdf7",
                                        X"c638",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"c638",
                                        X"c658",
                                        X"defb",
                                        X"ef7d",
                                        X"f7be",
                                        X"f7be",
                                        X"e0e4",
                                        X"e0e4",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"df7d",
                                        X"cf1c",
                                        X"cf1c",
                                        X"df5d",
                                        X"e0e4",
                                        X"df9e",
                                        X"efbe",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"d73d",
                                        X"c6dc",
                                        X"bedd",
                                        X"be7b",
                                        X"bdf8",
                                        X"bdf7",
                                        X"bdf8",
                                        X"be59",
                                        X"d71a",
                                        X"d75b",
                                        X"d75c",
                                        X"cf3c",
                                        X"bedc",
                                        X"be9b",
                                        X"bebc",
                                        X"be7b",
                                        X"be9b",
                                        X"bebc",
                                        X"be9b",
                                        X"c6bb",
                                        X"df3c",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef7d",
                                        X"e75c",
                                        X"e73c",
                                        X"defb",
                                        X"d6da",
                                        X"d6ba",
                                        X"ce99",
                                        X"d6ba",
                                        X"d6da",
                                        X"d6da",
                                        X"d69a",
                                        X"ce79",
                                        X"d69a",
                                        X"d6ba",
                                        X"d69a",
                                        X"d6da",
                                        X"e73c",
                                        X"ef7d",
                                        X"f7be",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"ef5c",
                                        X"d6ba",
                                        X"ef7d",
                                        X"e0e4",
                                        X"ef7d",
                                        X"d6da",
                                        X"e0e4",
                                        X"d6da",
                                        X"ce99",
                                        X"d6ba",
                                        X"d6ba",
                                        X"e0e4",
                                        X"ce79",
                                        X"ce99",
                                        X"e0e4",
                                        X"c658",
                                        X"be18",
                                        X"c638",
                                        X"e0e4",
                                        X"d6da",
                                        X"e73c",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"e0e4",
                                        X"e0e4",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"e0e4",
                                        X"d73d",
                                        X"cefc",
                                        X"d73d",
                                        X"e0e4",
                                        X"efde",
                                        X"f7de",
                                        X"e0e4",
                                        X"f7de",
                                        X"e7be",
                                        X"cf5e",
                                        X"e0e4",
                                        X"d75e",
                                        X"cf3e",
                                        X"c6db",
                                        X"c69a",
                                        X"c679",
                                        X"ced9",
                                        X"cf1a",
                                        X"d73b",
                                        X"d75b",
                                        X"cf3c",
                                        X"c6fc",
                                        X"c71c",
                                        X"bedc",
                                        X"bebc",
                                        X"be7b",
                                        X"bebc",
                                        X"bebb",
                                        X"be9a",
                                        X"cedb",
                                        X"e75d",
                                        X"ef9e",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef7d",
                                        X"e75c",
                                        X"e73c",
                                        X"defb",
                                        X"d6ba",
                                        X"d69a",
                                        X"d69a",
                                        X"d6da",
                                        X"d6da",
                                        X"df1b",
                                        X"d6da",
                                        X"d6ba",
                                        X"ce9a",
                                        X"d6ba",
                                        X"d6ba",
                                        X"d6da",
                                        X"e75c",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"f7de",
                                        X"f7be",
                                        X"df1b",
                                        X"e0e4",
                                        X"ef9d",
                                        X"ef7d",
                                        X"e0e4",
                                        X"c638",
                                        X"d6ba",
                                        X"defb",
                                        X"df1b",
                                        X"e0e4",
                                        X"ce79",
                                        X"ce59",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"ce99",
                                        X"e75d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7de",
                                        X"e0e4",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"f7de",
                                        X"e0e4",
                                        X"cefc",
                                        X"d73d",
                                        X"e0e4",
                                        X"d77e",
                                        X"e7be",
                                        X"e0e4",
                                        X"df9e",
                                        X"cf5e",
                                        X"cf5e",
                                        X"e0e4",
                                        X"df7e",
                                        X"df5c",
                                        X"d73b",
                                        X"cf1b",
                                        X"cf1a",
                                        X"d739",
                                        X"df59",
                                        X"d75b",
                                        X"df7c",
                                        X"d75c",
                                        X"bedc",
                                        X"c6fd",
                                        X"c6fd",
                                        X"bedd",
                                        X"bebc",
                                        X"be9b",
                                        X"be7a",
                                        X"be7a",
                                        X"cedc",
                                        X"ef7d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef7d",
                                        X"e75c",
                                        X"df1b",
                                        X"d6da",
                                        X"d6ba",
                                        X"d6da",
                                        X"d6da",
                                        X"defb",
                                        X"d6da",
                                        X"defb",
                                        X"ef7d",
                                        X"e75c",
                                        X"df1b",
                                        X"e73c",
                                        X"defb",
                                        X"defb",
                                        X"e75d",
                                        X"ef9e",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"e73c",
                                        X"e73c",
                                        X"e0e4",
                                        X"ce59",
                                        X"c638",
                                        X"ce59",
                                        X"c658",
                                        X"e0e4",
                                        X"ce79",
                                        X"ce79",
                                        X"e0e4",
                                        X"ef7d",
                                        X"e0e4",
                                        X"d6da",
                                        X"c658",
                                        X"d6da",
                                        X"ef7d",
                                        X"ef9d",
                                        X"f7be",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"f7de",
                                        X"ef9e",
                                        X"e0e4",
                                        X"c71d",
                                        X"e0e4",
                                        X"c73e",
                                        X"c75e",
                                        X"e0e4",
                                        X"cf7e",
                                        X"cf7e",
                                        X"cf5e",
                                        X"e0e4",
                                        X"df9d",
                                        X"d75c",
                                        X"df7c",
                                        X"df7a",
                                        X"d75a",
                                        X"d75a",
                                        X"d75a",
                                        X"df7c",
                                        X"df7c",
                                        X"cf5c",
                                        X"bedc",
                                        X"bebc",
                                        X"bedd",
                                        X"bedc",
                                        X"bebc",
                                        X"be9b",
                                        X"be9b",
                                        X"c69b",
                                        X"df1c",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"df1c",
                                        X"defb",
                                        X"d6da",
                                        X"d6da",
                                        X"d6da",
                                        X"defb",
                                        X"d6da",
                                        X"e73c",
                                        X"f7de",
                                        X"ef7d",
                                        X"ef9d",
                                        X"e75c",
                                        X"e73c",
                                        X"df1b",
                                        X"e75d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"ef7d",
                                        X"d6da",
                                        X"e0e4",
                                        X"d6ba",
                                        X"d6ba",
                                        X"c638",
                                        X"c638",
                                        X"e0e4",
                                        X"c658",
                                        X"d6db",
                                        X"e0e4",
                                        X"f7de",
                                        X"e75c",
                                        X"e0e4",
                                        X"ce59",
                                        X"c638",
                                        X"defb",
                                        X"ef7d",
                                        X"e0e4",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"f7de",
                                        X"f7de",
                                        X"df3d",
                                        X"e0e4",
                                        X"e0e4",
                                        X"bf3e",
                                        X"bf3e",
                                        X"e0e4",
                                        X"cf7e",
                                        X"cf5e",
                                        X"c73e",
                                        X"e0e4",
                                        X"cf3c",
                                        X"cf3c",
                                        X"df9c",
                                        X"d77a",
                                        X"d75b",
                                        X"d75c",
                                        X"d75c",
                                        X"cf3c",
                                        X"d73d",
                                        X"c6fc",
                                        X"befc",
                                        X"bedc",
                                        X"befd",
                                        X"bedd",
                                        X"bebb",
                                        X"be9b",
                                        X"be7a",
                                        X"cedb",
                                        X"e75d",
                                        X"efbe",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef7d",
                                        X"e75c",
                                        X"df1b",
                                        X"d6da",
                                        X"d6ba",
                                        X"d6ba",
                                        X"d6ba",
                                        X"d6da",
                                        X"d6da",
                                        X"e75c",
                                        X"f7de",
                                        X"e73c",
                                        X"df1c",
                                        X"e75c",
                                        X"e73c",
                                        X"df1b",
                                        X"ef7d",
                                        X"ef9d",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"ef9d",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"df1b",
                                        X"defb",
                                        X"e75c",
                                        X"ef7d",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"df1b",
                                        X"defb",
                                        X"e75c",
                                        X"e0e4",
                                        X"df1b",
                                        X"df1b",
                                        X"defb",
                                        X"e0e4",
                                        X"ce79",
                                        X"d6ba",
                                        X"ef7d",
                                        X"e0e4",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"f7de",
                                        X"f7de",
                                        X"e0e4",
                                        X"f7de",
                                        X"f7de",
                                        X"e77d",
                                        X"d71d",
                                        X"e0e4",
                                        X"bf1d",
                                        X"bf1d",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"e0e4",
                                        X"befd",
                                        X"bedc",
                                        X"cf1d",
                                        X"cf5c",
                                        X"cf3c",
                                        X"c71c",
                                        X"c6fd",
                                        X"c71d",
                                        X"bedc",
                                        X"cf3d",
                                        X"c6fc",
                                        X"bedc",
                                        X"c6fd",
                                        X"c6fd",
                                        X"bedd",
                                        X"be5a",
                                        X"be7a",
                                        X"be7a",
                                        X"d6fc",
                                        X"ef7d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"ef9d",
                                        X"e75d",
                                        X"e73c",
                                        X"defb",
                                        X"d6ba",
                                        X"d69a",
                                        X"d6ba",
                                        X"d6ba",
                                        X"d6da",
                                        X"df1b",
                                        X"e73c",
                                        X"e73c",
                                        X"f79e",
                                        X"e73c",
                                        X"d6ba",
                                        X"d69a",
                                        X"df1b",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"f7be",
                                        X"ef9d",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"ef7d",
                                        X"e75c",
                                        X"ef7d",
                                        X"e75c",
                                        X"defb",
                                        X"d6ba",
                                        X"ce79",
                                        X"df1b",
                                        X"e75c",
                                        X"defb",
                                        X"d6ba",
                                        X"d6ba",
                                        X"e73c",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e75d",
                                        X"c6fc",
                                        X"bedd",
                                        X"bf1d",
                                        X"bf3e",
                                        X"c75e",
                                        X"c73e",
                                        X"befd",
                                        X"bebc",
                                        X"bf1d",
                                        X"c71d",
                                        X"befd",
                                        X"c71d",
                                        X"befd",
                                        X"befd",
                                        X"c71d",
                                        X"bedd",
                                        X"c73e",
                                        X"c6fc",
                                        X"bebb",
                                        X"bedc",
                                        X"be9b",
                                        X"be9c",
                                        X"be5a",
                                        X"be5a",
                                        X"c6bb",
                                        X"e73c",
                                        X"ef9d",
                                        X"f7de",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"ef7d",
                                        X"e73c",
                                        X"e73c",
                                        X"defb",
                                        X"d6ba",
                                        X"ce79",
                                        X"ce99",
                                        X"d6ba",
                                        X"defb",
                                        X"df1b",
                                        X"e73c",
                                        X"e75c",
                                        X"e73c",
                                        X"d6ba",
                                        X"c658",
                                        X"ce79",
                                        X"e73c",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e75c",
                                        X"e75c",
                                        X"defb",
                                        X"e75c",
                                        X"e75c",
                                        X"e73c",
                                        X"e75c",
                                        X"d6da",
                                        X"d6da",
                                        X"df1c",
                                        X"ef9d",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"efbe",
                                        X"cedc",
                                        X"bedc",
                                        X"bf1e",
                                        X"befd",
                                        X"c73e",
                                        X"bf1d",
                                        X"be9c",
                                        X"befd",
                                        X"bf1e",
                                        X"bedd",
                                        X"befd",
                                        X"befd",
                                        X"befd",
                                        X"bf1e",
                                        X"befd",
                                        X"bedd",
                                        X"c71e",
                                        X"befd",
                                        X"bebc",
                                        X"bebc",
                                        X"be3a",
                                        X"be5a",
                                        X"be7a",
                                        X"be7a",
                                        X"d71c",
                                        X"ef7d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7be",
                                        X"f7be",
                                        X"ef7d",
                                        X"e75c",
                                        X"e73c",
                                        X"df1b",
                                        X"defb",
                                        X"d6ba",
                                        X"ce99",
                                        X"ce79",
                                        X"ce79",
                                        X"ce79",
                                        X"d6da",
                                        X"defb",
                                        X"ce99",
                                        X"c638",
                                        X"be17",
                                        X"c638",
                                        X"df1b",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7be",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"ef7d",
                                        X"e73c",
                                        X"ef7d",
                                        X"defb",
                                        X"d6da",
                                        X"df1b",
                                        X"e73c",
                                        X"e73c",
                                        X"defb",
                                        X"df1b",
                                        X"e75c",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e77d",
                                        X"bebc",
                                        X"befd",
                                        X"bedd",
                                        X"bedd",
                                        X"bedc",
                                        X"bedc",
                                        X"befd",
                                        X"bedd",
                                        X"be9c",
                                        X"befd",
                                        X"befd",
                                        X"befd",
                                        X"bedd",
                                        X"bedd",
                                        X"bedd",
                                        X"befd",
                                        X"bebc",
                                        X"be9b",
                                        X"be9c",
                                        X"be5b",
                                        X"be39",
                                        X"be7a",
                                        X"cedb",
                                        X"e75d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"ef9e",
                                        X"ef9d",
                                        X"ef7d",
                                        X"e75c",
                                        X"e75c",
                                        X"e73c",
                                        X"df1b",
                                        X"d6da",
                                        X"ce79",
                                        X"c638",
                                        X"c638",
                                        X"bdf7",
                                        X"bdf7",
                                        X"be17",
                                        X"c618",
                                        X"be18",
                                        X"c638",
                                        X"c658",
                                        X"d6ba",
                                        X"ef7d",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"ef7d",
                                        X"d6da",
                                        X"d6ba",
                                        X"e73c",
                                        X"e73c",
                                        X"d6da",
                                        X"e75c",
                                        X"e75c",
                                        X"defb",
                                        X"e75c",
                                        X"ef7d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"d73d",
                                        X"bebc",
                                        X"be9c",
                                        X"be9c",
                                        X"be9b",
                                        X"bebc",
                                        X"bedd",
                                        X"bedd",
                                        X"bebc",
                                        X"befd",
                                        X"bebc",
                                        X"bedc",
                                        X"bedd",
                                        X"bedd",
                                        X"bebc",
                                        X"bebc",
                                        X"be7b",
                                        X"be5a",
                                        X"be5a",
                                        X"be3a",
                                        X"be3a",
                                        X"c69b",
                                        X"df3c",
                                        X"ef9d",
                                        X"f79e",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e75c",
                                        X"e73c",
                                        X"defb",
                                        X"c658",
                                        X"c618",
                                        X"c618",
                                        X"c618",
                                        X"c638",
                                        X"c638",
                                        X"c618",
                                        X"c638",
                                        X"ce99",
                                        X"d6da",
                                        X"d6da",
                                        X"e75c",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"defb",
                                        X"d6da",
                                        X"e73c",
                                        X"e75c",
                                        X"ce99",
                                        X"df1b",
                                        X"e73c",
                                        X"ef7d",
                                        X"e75c",
                                        X"defb",
                                        X"e75c",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"d71c",
                                        X"be9b",
                                        X"be5a",
                                        X"be7b",
                                        X"be9c",
                                        X"bedd",
                                        X"bebc",
                                        X"be9c",
                                        X"bedd",
                                        X"be7b",
                                        X"be7b",
                                        X"bebc",
                                        X"be9c",
                                        X"be7b",
                                        X"be9c",
                                        X"be3a",
                                        X"be19",
                                        X"be39",
                                        X"be19",
                                        X"be7a",
                                        X"d6fb",
                                        X"e77d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e73c",
                                        X"df1c",
                                        X"defb",
                                        X"ce9a",
                                        X"c659",
                                        X"c658",
                                        X"c638",
                                        X"c618",
                                        X"be17",
                                        X"c638",
                                        X"c658",
                                        X"d6da",
                                        X"defb",
                                        X"e73c",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"d6da",
                                        X"df1b",
                                        X"e73c",
                                        X"ef7d",
                                        X"defb",
                                        X"e75c",
                                        X"e75c",
                                        X"defb",
                                        X"d6da",
                                        X"e73c",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"df3c",
                                        X"be9b",
                                        X"be9b",
                                        X"be7b",
                                        X"bebc",
                                        X"be5a",
                                        X"be5a",
                                        X"be9c",
                                        X"be5a",
                                        X"be5a",
                                        X"be5a",
                                        X"be5a",
                                        X"be7a",
                                        X"be5b",
                                        X"be39",
                                        X"be18",
                                        X"be39",
                                        X"be7a",
                                        X"d6fb",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"e75c",
                                        X"e73c",
                                        X"d6da",
                                        X"ce79",
                                        X"c638",
                                        X"be17",
                                        X"c638",
                                        X"c638",
                                        X"c638",
                                        X"c638",
                                        X"c658",
                                        X"ce79",
                                        X"ce59",
                                        X"defb",
                                        X"ef7d",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef9d",
                                        X"e73c",
                                        X"e75c",
                                        X"e75c",
                                        X"ef7d",
                                        X"df1b",
                                        X"d6da",
                                        X"e73c",
                                        X"df1b",
                                        X"df1b",
                                        X"e75c",
                                        X"d6db",
                                        X"e73c",
                                        X"ef7d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"e75d",
                                        X"cefb",
                                        X"be9a",
                                        X"be9b",
                                        X"be5a",
                                        X"be39",
                                        X"be5a",
                                        X"be5a",
                                        X"be39",
                                        X"be39",
                                        X"be39",
                                        X"be5a",
                                        X"be39",
                                        X"be39",
                                        X"be5a",
                                        X"c6bb",
                                        X"d71c",
                                        X"e75d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e75c",
                                        X"e73c",
                                        X"defb",
                                        X"d69a",
                                        X"c638",
                                        X"bdf7",
                                        X"be17",
                                        X"c658",
                                        X"ce79",
                                        X"c659",
                                        X"d6ba",
                                        X"d6ba",
                                        X"defb",
                                        X"defb",
                                        X"d6da",
                                        X"e73c",
                                        X"ef7d",
                                        X"ef7d",
                                        X"f7be",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"f7be",
                                        X"ef9d",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"defb",
                                        X"defb",
                                        X"e73c",
                                        X"e75c",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"e73c",
                                        X"defb",
                                        X"df1b",
                                        X"ef7d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"ef9d",
                                        X"e73c",
                                        X"d71c",
                                        X"cedb",
                                        X"be7a",
                                        X"be59",
                                        X"be5a",
                                        X"be5a",
                                        X"be5a",
                                        X"be5a",
                                        X"be5a",
                                        X"c67a",
                                        X"c69a",
                                        X"d6fb",
                                        X"e73c",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e75c",
                                        X"defb",
                                        X"defb",
                                        X"ce9a",
                                        X"c638",
                                        X"c659",
                                        X"c658",
                                        X"c658",
                                        X"c658",
                                        X"d6ba",
                                        X"d6db",
                                        X"d6da",
                                        X"df1b",
                                        X"df1b",
                                        X"e73c",
                                        X"e73c",
                                        X"e75c",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"f7de",
                                        X"e75c",
                                        X"d69a",
                                        X"d6da",
                                        X"d6da",
                                        X"e75c",
                                        X"defb",
                                        X"e75c",
                                        X"e73c",
                                        X"d6ba",
                                        X"ce59",
                                        X"d6ba",
                                        X"e73c",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"ef9d",
                                        X"e75d",
                                        X"df3c",
                                        X"d6fb",
                                        X"d6fb",
                                        X"d6db",
                                        X"d6db",
                                        X"d6db",
                                        X"d6fb",
                                        X"df1c",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e75d",
                                        X"e73c",
                                        X"defb",
                                        X"d6da",
                                        X"ce79",
                                        X"c638",
                                        X"ce79",
                                        X"d6ba",
                                        X"ce99",
                                        X"ce79",
                                        X"ce79",
                                        X"d6ba",
                                        X"d6da",
                                        X"d6da",
                                        X"e73c",
                                        X"e73c",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"f7be",
                                        X"f7be",
                                        X"ef9e",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ce99",
                                        X"d6ba",
                                        X"ce99",
                                        X"ce79",
                                        X"ce9a",
                                        X"ce79",
                                        X"ce59",
                                        X"ce9a",
                                        X"defb",
                                        X"e73c",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e75c",
                                        X"e73c",
                                        X"e73c",
                                        X"df1b",
                                        X"d6da",
                                        X"ce99",
                                        X"ce79",
                                        X"c658",
                                        X"ce79",
                                        X"ce99",
                                        X"c638",
                                        X"ce9a",
                                        X"d69a",
                                        X"d6ba",
                                        X"d6da",
                                        X"d6da",
                                        X"d6ba",
                                        X"df1b",
                                        X"e73c",
                                        X"e75c",
                                        X"e75c",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"ef7d",
                                        X"f7de",
                                        X"ef7d",
                                        X"f7be",
                                        X"ef9d",
                                        X"df1b",
                                        X"d6ba",
                                        X"ce79",
                                        X"ce99",
                                        X"ce99",
                                        X"d6da",
                                        X"ef7d",
                                        X"e75c",
                                        X"e73c",
                                        X"df1c",
                                        X"d69a",
                                        X"ce79",
                                        X"d6da",
                                        X"df1b",
                                        X"df1b",
                                        X"df1b",
                                        X"df1b",
                                        X"e71c",
                                        X"e73c",
                                        X"e73c",
                                        X"df1b",
                                        X"e75c",
                                        X"df1b",
                                        X"defb",
                                        X"defb",
                                        X"defb",
                                        X"defb",
                                        X"d6ba",
                                        X"d6ba",
                                        X"d6ba",
                                        X"d6ba",
                                        X"d6ba",
                                        X"d69a",
                                        X"d6da",
                                        X"defb",
                                        X"c658",
                                        X"d6da",
                                        X"defb",
                                        X"defb",
                                        X"ce99",
                                        X"ce99",
                                        X"ce79",
                                        X"d69a",
                                        X"defb",
                                        X"df1b",
                                        X"defb",
                                        X"df1b",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef9d",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9e",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"f79d",
                                        X"f79d",
                                        X"f7be",
                                        X"defb",
                                        X"d6da",
                                        X"df1b",
                                        X"defb",
                                        X"f7be",
                                        X"e75c",
                                        X"d6ba",
                                        X"dedb",
                                        X"defb",
                                        X"e73c",
                                        X"e75c",
                                        X"e75c",
                                        X"defb",
                                        X"d6ba",
                                        X"d6ba",
                                        X"ce79",
                                        X"d6ba",
                                        X"d6da",
                                        X"d6ba",
                                        X"ce9a",
                                        X"d6ba",
                                        X"d6ba",
                                        X"d69a",
                                        X"ce99",
                                        X"d6ba",
                                        X"c658",
                                        X"d69a",
                                        X"ce79",
                                        X"ce99",
                                        X"e73c",
                                        X"d6da",
                                        X"e73c",
                                        X"e75c",
                                        X"f7be",
                                        X"df1b",
                                        X"ce79",
                                        X"d6da",
                                        X"ce99",
                                        X"df1b",
                                        X"d6da",
                                        X"d6ba",
                                        X"d6ba",
                                        X"d6ba",
                                        X"df1c",
                                        X"df1b",
                                        X"e75c",
                                        X"e75c",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"d6da",
                                        X"e75c",
                                        X"e73c",
                                        X"f7de",
                                        X"e75c",
                                        X"ce99",
                                        X"ce79",
                                        X"d69a",
                                        X"d6ba",
                                        X"d6ba",
                                        X"d6da",
                                        X"ce99",
                                        X"ce99",
                                        X"df1b",
                                        X"defb",
                                        X"ce99",
                                        X"d6da",
                                        X"d6da",
                                        X"defb",
                                        X"e75c",
                                        X"e73c",
                                        X"defb",
                                        X"df1b",
                                        X"d6da",
                                        X"defb",
                                        X"d6ba",
                                        X"d6db",
                                        X"df1b",
                                        X"d6ba",
                                        X"d6da",
                                        X"d6ba",
                                        X"e73c",
                                        X"d6da",
                                        X"ef7d",
                                        X"defb",
                                        X"ce79",
                                        X"ce79",
                                        X"d69a",
                                        X"d69a",
                                        X"d6ba",
                                        X"d6da",
                                        X"defb",
                                        X"d6da",
                                        X"e73c",
                                        X"e73c",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9e",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"e75c",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef9d",
                                        X"e73c",
                                        X"df1b",
                                        X"e75c",
                                        X"ef7d",
                                        X"e73c",
                                        X"df1b",
                                        X"ef7d",
                                        X"d6da",
                                        X"ce99",
                                        X"e75c",
                                        X"df1b",
                                        X"e75c",
                                        X"d6db",
                                        X"ce99",
                                        X"defb",
                                        X"e75c",
                                        X"e73c",
                                        X"d6da",
                                        X"e73c",
                                        X"d6db",
                                        X"d6da",
                                        X"df1b",
                                        X"ef9d",
                                        X"d6ba",
                                        X"e73c",
                                        X"d6da",
                                        X"c659",
                                        X"ce99",
                                        X"ce99",
                                        X"d69a",
                                        X"defb",
                                        X"d6da",
                                        X"ce79",
                                        X"d69a",
                                        X"d6ba",
                                        X"d6da",
                                        X"d6da",
                                        X"d6da",
                                        X"defb",
                                        X"defb",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e75c",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"f79d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"ef7d",
                                        X"f7be",
                                        X"e75c",
                                        X"e73c",
                                        X"df1b",
                                        X"f7de",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"defb",
                                        X"d69a",
                                        X"ef9d",
                                        X"f79e",
                                        X"df1b",
                                        X"d6da",
                                        X"ce79",
                                        X"defb",
                                        X"d6db",
                                        X"ef7d",
                                        X"d6da",
                                        X"ce79",
                                        X"d6ba",
                                        X"e73c",
                                        X"defb",
                                        X"ce9a",
                                        X"e75c",
                                        X"df1b",
                                        X"d6ba",
                                        X"d6ba",
                                        X"d6ba",
                                        X"ce79",
                                        X"d6ba",
                                        X"d6ba",
                                        X"d6da",
                                        X"d6ba",
                                        X"ce99",
                                        X"d6ba",
                                        X"defb",
                                        X"df1b",
                                        X"defb",
                                        X"df1b",
                                        X"e75c",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"f7be",
                                        X"e73c",
                                        X"ef7d",
                                        X"f7de",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"ef9d",
                                        X"d6db",
                                        X"e73c",
                                        X"ef7d",
                                        X"e73c",
                                        X"ce9a",
                                        X"d6ba",
                                        X"df1b",
                                        X"e73c",
                                        X"df1b",
                                        X"e75d",
                                        X"d6ba",
                                        X"defb",
                                        X"d6da",
                                        X"d6da",
                                        X"ce79",
                                        X"defb",
                                        X"df1b",
                                        X"d6ba",
                                        X"ce79",
                                        X"d6ba",
                                        X"ce79",
                                        X"d6ba",
                                        X"d6da",
                                        X"ce99",
                                        X"d6ba",
                                        X"d6ba",
                                        X"d6ba",
                                        X"d6da",
                                        X"df1b",
                                        X"df1b",
                                        X"e73c",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e75c",
                                        X"ef7d",
                                        X"e75d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e75c",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"f7de",
                                        X"ef7d",
                                        X"f7bd",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"f7de",
                                        X"ef7d",
                                        X"defb",
                                        X"e75c",
                                        X"f7be",
                                        X"ef9d",
                                        X"e75c",
                                        X"defb",
                                        X"e75c",
                                        X"e73c",
                                        X"defb",
                                        X"df1b",
                                        X"e73c",
                                        X"d6da",
                                        X"defb",
                                        X"ce9a",
                                        X"ce99",
                                        X"d6da",
                                        X"ce99",
                                        X"ce79",
                                        X"d6ba",
                                        X"d6ba",
                                        X"d6ba",
                                        X"d6ba",
                                        X"d6da",
                                        X"ce99",
                                        X"d6ba",
                                        X"defb",
                                        X"d6da",
                                        X"defb",
                                        X"defb",
                                        X"e73c",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef9d",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"ef5c",
                                        X"ef7d",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e73c",
                                        X"defb",
                                        X"d6ba",
                                        X"d69a",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"d6da",
                                        X"d6ba",
                                        X"d6da",
                                        X"ce99",
                                        X"d6ba",
                                        X"d6da",
                                        X"defb",
                                        X"e73c",
                                        X"defb",
                                        X"e75c",
                                        X"e75c",
                                        X"ef9d",
                                        X"ef9d",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"e011",
                                        X"e011",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"f7be",
                                        X"ef9d",
                                        X"e011",
                                        X"ef9d",
                                        X"f7de",
                                        X"ef9d",
                                        X"f7be",
                                        X"e011",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"e011",
                                        X"d6da",
                                        X"d6ba",
                                        X"d6ba",
                                        X"e011",
                                        X"e73c",
                                        X"df1b",
                                        X"d6da",
                                        X"e011",
                                        X"d6ba",
                                        X"d6ba",
                                        X"d6db",
                                        X"df1b",
                                        X"e73c",
                                        X"e73c",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"e75c",
                                        X"e011",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e73c",
                                        X"e011",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e011",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e011",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"f7be",
                                        X"ef9d",
                                        X"e011",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"ef7d",
                                        X"e73c",
                                        X"df1b",
                                        X"defb",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e73c",
                                        X"df1c",
                                        X"e73c",
                                        X"e75c",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e75c",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e75c",
                                        X"e011",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e011",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"e011",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"ef9d",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"ef7d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7be",
                                        X"e011",
                                        X"f7de",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"e011",
                                        X"ef7d",
                                        X"e011",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"e73c",
                                        X"e75c",
                                        X"e011",
                                        X"e75c",
                                        X"e75c",
                                        X"e75c",
                                        X"e011",
                                        X"e75c",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef9d",
                                        X"e75d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e011",
                                        X"e011",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e011",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"ef9d",
                                        X"f7de",
                                        X"f7de",
                                        X"ef9d",
                                        X"e011",
                                        X"f7de",
                                        X"f79d",
                                        X"f7de",
                                        X"f7be",
                                        X"e011",
                                        X"ef7d",
                                        X"ef9e",
                                        X"e011",
                                        X"ef9d",
                                        X"e75c",
                                        X"e73c",
                                        X"e75c",
                                        X"e011",
                                        X"e75c",
                                        X"ef9d",
                                        X"f7be",
                                        X"e011",
                                        X"ef9d",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e011",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"e011",
                                        X"f79e",
                                        X"f7be",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"f7de",
                                        X"f79d",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"f7de",
                                        X"f7be",
                                        X"e011",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"e011",
                                        X"ef7d",
                                        X"e73c",
                                        X"ef9d",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"ef9d",
                                        X"f79e",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9e",
                                        X"f7be",
                                        X"e011",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"e011",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"e011",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f79d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7be",
                                        X"f7be",
                                        X"ef9d",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"ef9e",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"f7de",
                                        X"f7be",
                                        X"f7de",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9e",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"ef9e",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef7d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7be",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f483",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7be",
                                        X"f7be",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"ef9d",
                                        X"f7be",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de",
                                        X"f7de"
                                    );
    signal sdata_out1   : STD_LOGIC_VECTOR (15 downto 0);
    signal sdata_out2   : STD_LOGIC_VECTOR (15 downto 0);
    
begin

    process(address1, mem)
        begin
            sdata_out1 <= mem(to_integer(unsigned(address1)));
    end process;
    
    data_out1   <= sdata_out1;
    
    process(address2, mem)
        begin
            sdata_out2 <= mem(to_integer(unsigned(address2)));
    end process;
    
    data_out2   <= sdata_out2;
    
    process(clk1, reset)
        begin
            if rising_edge(clk1) then
                if w2 = '1' then
                    mem(to_integer(unsigned(address2))) <= data_in2;
                end if;
            end if;
    end process;
    
end Behavioral;